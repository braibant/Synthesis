// tag associated with this file
//adder4_0.1
module Adder (clk, rst_n, guard, value, reg_0, reg_1);
integer index; // Used for initialisations
input clk;
input rst_n;
output guard;
output [33:0] value;
// state declarations
input [15:0] reg_0;
input [15:0] reg_1;
// bindings 
wire  wire0 = 0'b0;
wire  wire1 = 1'b1;
wire  wire2 = 1'b0;
wire [15:0] wire3 = reg_1;
wire [15:0] wire4 = reg_0;
wire [7:0] wire5 = wire3[7:0];
wire [7:0] wire6 = wire3[15:8];
wire [7:0] wire7 = wire4[7:0];
wire [7:0] wire8 = wire4[15:8];
wire [3:0] wire9 = wire5[3:0];
wire [3:0] wire10 = wire5[7:4];
wire [3:0] wire11 = wire7[3:0];
wire [3:0] wire12 = wire7[7:4];
wire [1:0] wire13 = wire9[1:0];
wire [1:0] wire14 = wire9[3:2];
wire [1:0] wire15 = wire11[1:0];
wire [1:0] wire16 = wire11[3:2];
wire  wire17 = wire13[0:0];
wire  wire18 = wire13[1:1];
wire  wire19 = wire15[0:0];
wire  wire20 = wire15[1:1];
wire  wire21 = 1'b1;
wire  wire22 = wire17 == wire21;
wire  wire23 = wire19 == wire21;
wire  wire24 = wire22 | wire23;
wire  wire25 = wire22 & wire23;
wire  wire26 = wire17 + wire19;
wire  wire27 = wire26 + wire21;
wire [3:0] wire28 = {wire24, wire25, wire26, wire27};
wire  wire29 = wire18 == wire21;
wire  wire30 = wire20 == wire21;
wire  wire31 = wire29 | wire30;
wire  wire32 = wire29 & wire30;
wire  wire33 = wire18 + wire20;
wire  wire34 = wire33 + wire21;
wire [3:0] wire35 = {wire31, wire32, wire33, wire34};
wire [2:0] wire36 = wire28[3:1];
wire [1:0] wire37 = wire36[2:1];
wire  wire38 = wire37[1:1];
wire  wire39 = 0;
wire [2:0] wire40 = wire35[3:1];
wire [1:0] wire41 = wire40[2:1];
wire  wire42 = wire41[1:1];
wire  wire43 = wire25 ? wire34 : wire33;
wire  wire44 = wire24 ? wire34 : wire33;
wire  wire45 = wire31 & wire24;
wire  wire46 = wire32 | wire45;
wire  wire47 = wire31 & wire25;
wire  wire48 = wire32 | wire47;
wire [1:0] wire49 = {wire43, wire26};
wire [1:0] wire50 = {wire44, wire27};
wire [5:0] wire51 = {wire46, wire48, wire49, wire50};
wire  wire52 = wire14[0:0];
wire  wire53 = wire14[1:1];
wire  wire54 = wire16[0:0];
wire  wire55 = wire16[1:1];
wire  wire56 = wire52 == wire21;
wire  wire57 = wire54 == wire21;
wire  wire58 = wire56 | wire57;
wire  wire59 = wire56 & wire57;
wire  wire60 = wire52 + wire54;
wire  wire61 = wire60 + wire21;
wire [3:0] wire62 = {wire58, wire59, wire60, wire61};
wire  wire63 = wire53 == wire21;
wire  wire64 = wire55 == wire21;
wire  wire65 = wire63 | wire64;
wire  wire66 = wire63 & wire64;
wire  wire67 = wire53 + wire55;
wire  wire68 = wire67 + wire21;
wire [3:0] wire69 = {wire65, wire66, wire67, wire68};
wire [2:0] wire70 = wire62[3:1];
wire [1:0] wire71 = wire70[2:1];
wire  wire72 = wire71[1:1];
wire [2:0] wire73 = wire69[3:1];
wire [1:0] wire74 = wire73[2:1];
wire  wire75 = wire74[1:1];
wire  wire76 = wire59 ? wire68 : wire67;
wire  wire77 = wire58 ? wire68 : wire67;
wire  wire78 = wire65 & wire58;
wire  wire79 = wire66 | wire78;
wire  wire80 = wire65 & wire59;
wire  wire81 = wire66 | wire80;
wire [1:0] wire82 = {wire76, wire60};
wire [1:0] wire83 = {wire77, wire61};
wire [5:0] wire84 = {wire79, wire81, wire82, wire83};
wire [4:0] wire85 = wire51[5:1];
wire [3:0] wire86 = wire85[4:1];
wire [1:0] wire87 = wire86[3:2];
wire [4:0] wire88 = wire84[5:1];
wire [3:0] wire89 = wire88[4:1];
wire [1:0] wire90 = wire89[3:2];
wire [1:0] wire91 = wire48 ? wire83 : wire82;
wire [1:0] wire92 = wire46 ? wire83 : wire82;
wire  wire93 = wire79 & wire46;
wire  wire94 = wire81 | wire93;
wire  wire95 = wire79 & wire48;
wire  wire96 = wire81 | wire95;
wire [3:0] wire97 = {wire91, wire49};
wire [3:0] wire98 = {wire92, wire50};
wire [9:0] wire99 = {wire94, wire96, wire97, wire98};
wire [1:0] wire100 = wire10[1:0];
wire [1:0] wire101 = wire10[3:2];
wire [1:0] wire102 = wire12[1:0];
wire [1:0] wire103 = wire12[3:2];
wire  wire104 = wire100[0:0];
wire  wire105 = wire100[1:1];
wire  wire106 = wire102[0:0];
wire  wire107 = wire102[1:1];
wire  wire108 = wire104 == wire21;
wire  wire109 = wire106 == wire21;
wire  wire110 = wire108 | wire109;
wire  wire111 = wire108 & wire109;
wire  wire112 = wire104 + wire106;
wire  wire113 = wire112 + wire21;
wire [3:0] wire114 = {wire110, wire111, wire112, wire113};
wire  wire115 = wire105 == wire21;
wire  wire116 = wire107 == wire21;
wire  wire117 = wire115 | wire116;
wire  wire118 = wire115 & wire116;
wire  wire119 = wire105 + wire107;
wire  wire120 = wire119 + wire21;
wire [3:0] wire121 = {wire117, wire118, wire119, wire120};
wire [2:0] wire122 = wire114[3:1];
wire [1:0] wire123 = wire122[2:1];
wire  wire124 = wire123[1:1];
wire [2:0] wire125 = wire121[3:1];
wire [1:0] wire126 = wire125[2:1];
wire  wire127 = wire126[1:1];
wire  wire128 = wire111 ? wire120 : wire119;
wire  wire129 = wire110 ? wire120 : wire119;
wire  wire130 = wire117 & wire110;
wire  wire131 = wire118 | wire130;
wire  wire132 = wire117 & wire111;
wire  wire133 = wire118 | wire132;
wire [1:0] wire134 = {wire128, wire112};
wire [1:0] wire135 = {wire129, wire113};
wire [5:0] wire136 = {wire131, wire133, wire134, wire135};
wire  wire137 = wire101[0:0];
wire  wire138 = wire101[1:1];
wire  wire139 = wire103[0:0];
wire  wire140 = wire103[1:1];
wire  wire141 = wire137 == wire21;
wire  wire142 = wire139 == wire21;
wire  wire143 = wire141 | wire142;
wire  wire144 = wire141 & wire142;
wire  wire145 = wire137 + wire139;
wire  wire146 = wire145 + wire21;
wire [3:0] wire147 = {wire143, wire144, wire145, wire146};
wire  wire148 = wire138 == wire21;
wire  wire149 = wire140 == wire21;
wire  wire150 = wire148 | wire149;
wire  wire151 = wire148 & wire149;
wire  wire152 = wire138 + wire140;
wire  wire153 = wire152 + wire21;
wire [3:0] wire154 = {wire150, wire151, wire152, wire153};
wire [2:0] wire155 = wire147[3:1];
wire [1:0] wire156 = wire155[2:1];
wire  wire157 = wire156[1:1];
wire [2:0] wire158 = wire154[3:1];
wire [1:0] wire159 = wire158[2:1];
wire  wire160 = wire159[1:1];
wire  wire161 = wire144 ? wire153 : wire152;
wire  wire162 = wire143 ? wire153 : wire152;
wire  wire163 = wire150 & wire143;
wire  wire164 = wire151 | wire163;
wire  wire165 = wire150 & wire144;
wire  wire166 = wire151 | wire165;
wire [1:0] wire167 = {wire161, wire145};
wire [1:0] wire168 = {wire162, wire146};
wire [5:0] wire169 = {wire164, wire166, wire167, wire168};
wire [4:0] wire170 = wire136[5:1];
wire [3:0] wire171 = wire170[4:1];
wire [1:0] wire172 = wire171[3:2];
wire [4:0] wire173 = wire169[5:1];
wire [3:0] wire174 = wire173[4:1];
wire [1:0] wire175 = wire174[3:2];
wire [1:0] wire176 = wire133 ? wire168 : wire167;
wire [1:0] wire177 = wire131 ? wire168 : wire167;
wire  wire178 = wire164 & wire131;
wire  wire179 = wire166 | wire178;
wire  wire180 = wire164 & wire133;
wire  wire181 = wire166 | wire180;
wire [3:0] wire182 = {wire176, wire134};
wire [3:0] wire183 = {wire177, wire135};
wire [9:0] wire184 = {wire179, wire181, wire182, wire183};
wire [8:0] wire185 = wire99[9:1];
wire [7:0] wire186 = wire185[8:1];
wire [3:0] wire187 = wire186[7:4];
wire [8:0] wire188 = wire184[9:1];
wire [7:0] wire189 = wire188[8:1];
wire [3:0] wire190 = wire189[7:4];
wire [3:0] wire191 = wire96 ? wire183 : wire182;
wire [3:0] wire192 = wire94 ? wire183 : wire182;
wire  wire193 = wire179 & wire94;
wire  wire194 = wire181 | wire193;
wire  wire195 = wire179 & wire96;
wire  wire196 = wire181 | wire195;
wire [7:0] wire197 = {wire191, wire97};
wire [7:0] wire198 = {wire192, wire98};
wire [17:0] wire199 = {wire194, wire196, wire197, wire198};
wire [3:0] wire200 = wire6[3:0];
wire [3:0] wire201 = wire6[7:4];
wire [3:0] wire202 = wire8[3:0];
wire [3:0] wire203 = wire8[7:4];
wire [1:0] wire204 = wire200[1:0];
wire [1:0] wire205 = wire200[3:2];
wire [1:0] wire206 = wire202[1:0];
wire [1:0] wire207 = wire202[3:2];
wire  wire208 = wire204[0:0];
wire  wire209 = wire204[1:1];
wire  wire210 = wire206[0:0];
wire  wire211 = wire206[1:1];
wire  wire212 = wire208 == wire21;
wire  wire213 = wire210 == wire21;
wire  wire214 = wire212 | wire213;
wire  wire215 = wire212 & wire213;
wire  wire216 = wire208 + wire210;
wire  wire217 = wire216 + wire21;
wire [3:0] wire218 = {wire214, wire215, wire216, wire217};
wire  wire219 = wire209 == wire21;
wire  wire220 = wire211 == wire21;
wire  wire221 = wire219 | wire220;
wire  wire222 = wire219 & wire220;
wire  wire223 = wire209 + wire211;
wire  wire224 = wire223 + wire21;
wire [3:0] wire225 = {wire221, wire222, wire223, wire224};
wire [2:0] wire226 = wire218[3:1];
wire [1:0] wire227 = wire226[2:1];
wire  wire228 = wire227[1:1];
wire [2:0] wire229 = wire225[3:1];
wire [1:0] wire230 = wire229[2:1];
wire  wire231 = wire230[1:1];
wire  wire232 = wire215 ? wire224 : wire223;
wire  wire233 = wire214 ? wire224 : wire223;
wire  wire234 = wire221 & wire214;
wire  wire235 = wire222 | wire234;
wire  wire236 = wire221 & wire215;
wire  wire237 = wire222 | wire236;
wire [1:0] wire238 = {wire232, wire216};
wire [1:0] wire239 = {wire233, wire217};
wire [5:0] wire240 = {wire235, wire237, wire238, wire239};
wire  wire241 = wire205[0:0];
wire  wire242 = wire205[1:1];
wire  wire243 = wire207[0:0];
wire  wire244 = wire207[1:1];
wire  wire245 = wire241 == wire21;
wire  wire246 = wire243 == wire21;
wire  wire247 = wire245 | wire246;
wire  wire248 = wire245 & wire246;
wire  wire249 = wire241 + wire243;
wire  wire250 = wire249 + wire21;
wire [3:0] wire251 = {wire247, wire248, wire249, wire250};
wire  wire252 = wire242 == wire21;
wire  wire253 = wire244 == wire21;
wire  wire254 = wire252 | wire253;
wire  wire255 = wire252 & wire253;
wire  wire256 = wire242 + wire244;
wire  wire257 = wire256 + wire21;
wire [3:0] wire258 = {wire254, wire255, wire256, wire257};
wire [2:0] wire259 = wire251[3:1];
wire [1:0] wire260 = wire259[2:1];
wire  wire261 = wire260[1:1];
wire [2:0] wire262 = wire258[3:1];
wire [1:0] wire263 = wire262[2:1];
wire  wire264 = wire263[1:1];
wire  wire265 = wire248 ? wire257 : wire256;
wire  wire266 = wire247 ? wire257 : wire256;
wire  wire267 = wire254 & wire247;
wire  wire268 = wire255 | wire267;
wire  wire269 = wire254 & wire248;
wire  wire270 = wire255 | wire269;
wire [1:0] wire271 = {wire265, wire249};
wire [1:0] wire272 = {wire266, wire250};
wire [5:0] wire273 = {wire268, wire270, wire271, wire272};
wire [4:0] wire274 = wire240[5:1];
wire [3:0] wire275 = wire274[4:1];
wire [1:0] wire276 = wire275[3:2];
wire [4:0] wire277 = wire273[5:1];
wire [3:0] wire278 = wire277[4:1];
wire [1:0] wire279 = wire278[3:2];
wire [1:0] wire280 = wire237 ? wire272 : wire271;
wire [1:0] wire281 = wire235 ? wire272 : wire271;
wire  wire282 = wire268 & wire235;
wire  wire283 = wire270 | wire282;
wire  wire284 = wire268 & wire237;
wire  wire285 = wire270 | wire284;
wire [3:0] wire286 = {wire280, wire238};
wire [3:0] wire287 = {wire281, wire239};
wire [9:0] wire288 = {wire283, wire285, wire286, wire287};
wire [1:0] wire289 = wire201[1:0];
wire [1:0] wire290 = wire201[3:2];
wire [1:0] wire291 = wire203[1:0];
wire [1:0] wire292 = wire203[3:2];
wire  wire293 = wire289[0:0];
wire  wire294 = wire289[1:1];
wire  wire295 = wire291[0:0];
wire  wire296 = wire291[1:1];
wire  wire297 = wire293 == wire21;
wire  wire298 = wire295 == wire21;
wire  wire299 = wire297 | wire298;
wire  wire300 = wire297 & wire298;
wire  wire301 = wire293 + wire295;
wire  wire302 = wire301 + wire21;
wire [3:0] wire303 = {wire299, wire300, wire301, wire302};
wire  wire304 = wire294 == wire21;
wire  wire305 = wire296 == wire21;
wire  wire306 = wire304 | wire305;
wire  wire307 = wire304 & wire305;
wire  wire308 = wire294 + wire296;
wire  wire309 = wire308 + wire21;
wire [3:0] wire310 = {wire306, wire307, wire308, wire309};
wire [2:0] wire311 = wire303[3:1];
wire [1:0] wire312 = wire311[2:1];
wire  wire313 = wire312[1:1];
wire [2:0] wire314 = wire310[3:1];
wire [1:0] wire315 = wire314[2:1];
wire  wire316 = wire315[1:1];
wire  wire317 = wire300 ? wire309 : wire308;
wire  wire318 = wire299 ? wire309 : wire308;
wire  wire319 = wire306 & wire299;
wire  wire320 = wire307 | wire319;
wire  wire321 = wire306 & wire300;
wire  wire322 = wire307 | wire321;
wire [1:0] wire323 = {wire317, wire301};
wire [1:0] wire324 = {wire318, wire302};
wire [5:0] wire325 = {wire320, wire322, wire323, wire324};
wire  wire326 = wire290[0:0];
wire  wire327 = wire290[1:1];
wire  wire328 = wire292[0:0];
wire  wire329 = wire292[1:1];
wire  wire330 = wire326 == wire21;
wire  wire331 = wire328 == wire21;
wire  wire332 = wire330 | wire331;
wire  wire333 = wire330 & wire331;
wire  wire334 = wire326 + wire328;
wire  wire335 = wire334 + wire21;
wire [3:0] wire336 = {wire332, wire333, wire334, wire335};
wire  wire337 = wire327 == wire21;
wire  wire338 = wire329 == wire21;
wire  wire339 = wire337 | wire338;
wire  wire340 = wire337 & wire338;
wire  wire341 = wire327 + wire329;
wire  wire342 = wire341 + wire21;
wire [3:0] wire343 = {wire339, wire340, wire341, wire342};
wire [2:0] wire344 = wire336[3:1];
wire [1:0] wire345 = wire344[2:1];
wire  wire346 = wire345[1:1];
wire [2:0] wire347 = wire343[3:1];
wire [1:0] wire348 = wire347[2:1];
wire  wire349 = wire348[1:1];
wire  wire350 = wire333 ? wire342 : wire341;
wire  wire351 = wire332 ? wire342 : wire341;
wire  wire352 = wire339 & wire332;
wire  wire353 = wire340 | wire352;
wire  wire354 = wire339 & wire333;
wire  wire355 = wire340 | wire354;
wire [1:0] wire356 = {wire350, wire334};
wire [1:0] wire357 = {wire351, wire335};
wire [5:0] wire358 = {wire353, wire355, wire356, wire357};
wire [4:0] wire359 = wire325[5:1];
wire [3:0] wire360 = wire359[4:1];
wire [1:0] wire361 = wire360[3:2];
wire [4:0] wire362 = wire358[5:1];
wire [3:0] wire363 = wire362[4:1];
wire [1:0] wire364 = wire363[3:2];
wire [1:0] wire365 = wire322 ? wire357 : wire356;
wire [1:0] wire366 = wire320 ? wire357 : wire356;
wire  wire367 = wire353 & wire320;
wire  wire368 = wire355 | wire367;
wire  wire369 = wire353 & wire322;
wire  wire370 = wire355 | wire369;
wire [3:0] wire371 = {wire365, wire323};
wire [3:0] wire372 = {wire366, wire324};
wire [9:0] wire373 = {wire368, wire370, wire371, wire372};
wire [8:0] wire374 = wire288[9:1];
wire [7:0] wire375 = wire374[8:1];
wire [3:0] wire376 = wire375[7:4];
wire [8:0] wire377 = wire373[9:1];
wire [7:0] wire378 = wire377[8:1];
wire [3:0] wire379 = wire378[7:4];
wire [3:0] wire380 = wire285 ? wire372 : wire371;
wire [3:0] wire381 = wire283 ? wire372 : wire371;
wire  wire382 = wire368 & wire283;
wire  wire383 = wire370 | wire382;
wire  wire384 = wire368 & wire285;
wire  wire385 = wire370 | wire384;
wire [7:0] wire386 = {wire380, wire286};
wire [7:0] wire387 = {wire381, wire287};
wire [17:0] wire388 = {wire383, wire385, wire386, wire387};
wire [16:0] wire389 = wire199[17:1];
wire [15:0] wire390 = wire389[16:1];
wire [7:0] wire391 = wire390[15:8];
wire [16:0] wire392 = wire388[17:1];
wire [15:0] wire393 = wire392[16:1];
wire [7:0] wire394 = wire393[15:8];
wire [7:0] wire395 = wire196 ? wire387 : wire386;
wire [7:0] wire396 = wire194 ? wire387 : wire386;
wire  wire397 = wire383 & wire194;
wire  wire398 = wire385 | wire397;
wire  wire399 = wire383 & wire196;
wire  wire400 = wire385 | wire399;
wire [15:0] wire401 = {wire395, wire197};
wire [15:0] wire402 = {wire396, wire198};
wire [33:0] wire403 = {wire398, wire400, wire401, wire402};
// effects 
assign guard = wire1;
assign value = wire403;
always@(posedge clk)
begin
	if(rst_n)
		begin
// reset 
		end
	else
		begin
	if(wire1)
		begin
// put  debug code here (display, stop, ...)
		end
		end
end
endmodule
