module Stack (clk, rst_n, guard, value);
integer index; // Used for initialisations
input clk;
input rst_n;
output guard;
output [0:0] value;
// state declarations
reg [7:0] reg_0 [255:0];
reg [7:0] reg_1 [255:0];
reg [7:0] reg_2;
reg [11:0] reg_3 [255:0];
reg [7:0] reg_4;
// bindings 
wire  wire0 = 0'b0;
wire  wire1 = 1'b1;
wire  wire2 = 1'b0;
wire [7:0] wire3 = reg_4;
wire [11:0] wire4 = reg_3[wire3];
wire [3:0] wire5 = wire4[3:0];
wire [3:0] wire6 = 4'b0;
wire  wire7 = wire5 == wire6;
wire [7:0] wire8 = reg_2;
wire [7:0] wire9 = wire4[11:4];
wire [7:0] wire10 = 8'b1;
wire [7:0] wire11 = wire8 + wire10;
wire [7:0] wire12 = wire3 + wire10;
wire [11:0] wire13 = reg_3[wire3];
wire [3:0] wire14 = wire13[3:0];
wire [3:0] wire15 = 4'b1;
wire  wire16 = wire14 == wire15;
wire [7:0] wire17 = wire13[11:4];
wire [7:0] wire18 = reg_0[wire17];
wire [11:0] wire19 = reg_3[wire3];
wire [3:0] wire20 = wire19[3:0];
wire [3:0] wire21 = 4'b10;
wire  wire22 = wire20 == wire21;
wire [7:0] wire23 = wire8 - wire10;
wire [7:0] wire24 = reg_1[wire23];
wire [7:0] wire25 = wire19[11:4];
wire  wire26 = wire7 | wire16;
wire [11:0] wire27 = reg_3[wire3];
wire [3:0] wire28 = wire27[3:0];
wire [3:0] wire29 = 4'b11;
wire  wire30 = wire28 == wire29;
wire [7:0] wire31 = reg_1[wire23];
wire [7:0] wire32 = 8'b10;
wire [7:0] wire33 = wire8 - wire32;
wire [7:0] wire34 = reg_1[wire33];
wire [7:0] wire35 = wire34 + wire31;
wire  wire36 = wire26 | wire22;
wire [11:0] wire37 = reg_3[wire3];
wire [3:0] wire38 = wire37[3:0];
wire [3:0] wire39 = 4'b100;
wire  wire40 = wire38 == wire39;
wire [7:0] wire41 = reg_1[wire23];
wire [7:0] wire42 = reg_1[wire33];
wire [7:0] wire43 = wire42 - wire41;
wire  wire44 = wire36 | wire30;
wire [11:0] wire45 = reg_3[wire3];
wire [3:0] wire46 = wire45[3:0];
wire [3:0] wire47 = 4'b101;
wire  wire48 = wire46 == wire47;
wire [7:0] wire49 = wire45[11:4];
wire [7:0] wire50 = wire12 + wire49;
wire  wire51 = wire44 | wire40;
wire [11:0] wire52 = reg_3[wire3];
wire [3:0] wire53 = wire52[3:0];
wire [3:0] wire54 = 4'b110;
wire  wire55 = wire53 == wire54;
wire [7:0] wire56 = wire52[11:4];
wire [7:0] wire57 = wire12 - wire56;
wire  wire58 = wire51 | wire48;
wire [11:0] wire59 = reg_3[wire3];
wire [3:0] wire60 = wire59[3:0];
wire [3:0] wire61 = 4'b111;
wire  wire62 = wire60 == wire61;
wire [7:0] wire63 = reg_1[wire23];
wire [7:0] wire64 = reg_1[wire33];
wire  wire65 = wire64 == wire63;
wire [7:0] wire66 = wire59[11:4];
wire [7:0] wire67 = wire12 + wire66;
wire  wire68 = wire58 | wire55;
wire [11:0] wire69 = reg_3[wire3];
wire [3:0] wire70 = wire69[3:0];
wire [3:0] wire71 = 4'b1001;
wire  wire72 = wire70 == wire71;
wire [7:0] wire73 = reg_1[wire23];
wire [7:0] wire74 = reg_1[wire33];
wire  wire75 = wire74 < wire73;
wire  wire76 = wire74 == wire73;
wire  wire77 = wire75 | wire76;
wire [7:0] wire78 = wire69[11:4];
wire [7:0] wire79 = wire12 + wire78;
wire  wire80 = wire68 | wire62;
wire [11:0] wire81 = reg_3[wire3];
wire [3:0] wire82 = wire81[3:0];
wire [3:0] wire83 = 4'b1010;
wire  wire84 = wire82 == wire83;
wire [7:0] wire85 = reg_1[wire23];
wire [7:0] wire86 = reg_1[wire33];
wire  wire87 = wire85 < wire86;
wire [7:0] wire88 = wire81[11:4];
wire [7:0] wire89 = wire12 + wire88;
wire  wire90 = wire80 | wire72;
wire [11:0] wire91 = reg_3[wire3];
wire [3:0] wire92 = wire91[3:0];
wire [3:0] wire93 = 4'b1011;
wire  wire94 = wire92 == wire93;
wire  wire95 = wire90 | wire84;
wire  wire96 = wire95 ? wire2 : wire1;
wire  wire97 = wire95 | wire94;
wire  wire98 = wire26 & wire7;
wire  wire99 = ~ wire7;
wire  wire100 = wire99 & wire16;
wire [7:0] wire101 = wire98 ? wire9 : wire18;
wire  wire102 = ~ wire26;
wire  wire103 = wire102 & wire22;
wire [7:0] wire104 = wire26 ? wire11 : wire23;
wire  wire105 = ~ wire36;
wire  wire106 = wire105 & wire30;
wire  wire107 = wire26 | wire106;
wire [7:0] wire108 = wire26 ? wire8 : wire33;
wire [7:0] wire109 = wire26 ? wire101 : wire35;
wire [7:0] wire110 = wire36 ? wire104 : wire23;
wire  wire111 = ~ wire44;
wire  wire112 = wire111 & wire40;
wire  wire113 = wire107 | wire112;
wire [7:0] wire114 = wire107 ? wire108 : wire33;
wire [7:0] wire115 = wire107 ? wire109 : wire43;
wire [7:0] wire116 = wire44 ? wire110 : wire23;
wire  wire117 = ~ wire51;
wire  wire118 = wire117 & wire48;
wire [7:0] wire119 = wire51 ? wire12 : wire50;
wire  wire120 = ~ wire58;
wire  wire121 = wire120 & wire55;
wire [7:0] wire122 = wire58 ? wire119 : wire57;
wire  wire123 = ~ wire68;
wire  wire124 = wire123 & wire62;
wire  wire125 = wire51 | wire124;
wire [7:0] wire126 = wire51 ? wire116 : wire33;
wire  wire127 = wire124 & wire65;
wire  wire128 = wire68 | wire127;
wire [7:0] wire129 = wire68 ? wire122 : wire67;
wire  wire130 = ~ wire65;
wire  wire131 = wire124 & wire130;
wire [7:0] wire132 = wire128 ? wire129 : wire12;
wire  wire133 = ~ wire80;
wire  wire134 = wire133 & wire72;
wire  wire135 = wire125 | wire134;
wire [7:0] wire136 = wire125 ? wire126 : wire33;
wire  wire137 = wire134 & wire77;
wire  wire138 = wire80 | wire137;
wire [7:0] wire139 = wire80 ? wire132 : wire79;
wire  wire140 = ~ wire77;
wire  wire141 = wire134 & wire140;
wire [7:0] wire142 = wire138 ? wire139 : wire12;
wire  wire143 = ~ wire90;
wire  wire144 = wire143 & wire84;
wire  wire145 = wire135 | wire144;
wire [7:0] wire146 = wire135 ? wire136 : wire33;
wire  wire147 = wire144 & wire87;
wire  wire148 = wire90 | wire147;
wire [7:0] wire149 = wire90 ? wire142 : wire89;
wire  wire150 = ~ wire87;
wire  wire151 = wire144 & wire150;
wire [7:0] wire152 = wire148 ? wire149 : wire12;
// effects 
assign guard = wire97;
assign value = wire96;
always@(posedge clk)
begin
	if(rst_n)
		begin
// reset 
		end
	else
		begin
// put  debug code here (display, stop, ...)
if(wire95) reg_4 <= wire152;
if(wire145) reg_2 <= wire146;
if(wire113) reg_1[wire114] <= wire115;
if(wire103) reg_0[wire25] <= wire24;
		end
end
endmodule
