module Sorter (clk, rst_n, guard, value, reg_0);
integer index; // Used for initialisations
input clk;
input rst_n;
output guard;
output [63:0] value;
// state declarations
input [63:0] reg_0;
// bindings 
wire  wire0 = 0'b0;
wire  wire1 = 1'b1;
wire  wire2 = 1'b0;
wire [63:0] wire3 = reg_0;
wire [31:0] wire4 = wire3[31:0];
wire [31:0] wire5 = wire3[63:32];
wire [31:0] wire6 = wire5[31:0];
wire [15:0] wire7 = wire4[15:0];
wire [15:0] wire8 = wire4[31:16];
wire [15:0] wire9 = wire8[15:0];
wire [7:0] wire10 = wire7[7:0];
wire [7:0] wire11 = wire7[15:8];
wire [7:0] wire12 = wire11[7:0];
wire [3:0] wire13 = wire10[3:0];
wire [3:0] wire14 = wire10[7:4];
wire [3:0] wire15 = wire14[3:0];
wire [3:0] wire16 = wire12[3:0];
wire [3:0] wire17 = wire12[7:4];
wire [3:0] wire18 = wire17[3:0];
wire [7:0] wire19 = wire9[7:0];
wire [7:0] wire20 = wire9[15:8];
wire [7:0] wire21 = wire20[7:0];
wire [3:0] wire22 = wire19[3:0];
wire [3:0] wire23 = wire19[7:4];
wire [3:0] wire24 = wire23[3:0];
wire [3:0] wire25 = wire21[3:0];
wire [3:0] wire26 = wire21[7:4];
wire [3:0] wire27 = wire26[3:0];
wire [15:0] wire28 = wire6[15:0];
wire [15:0] wire29 = wire6[31:16];
wire [15:0] wire30 = wire29[15:0];
wire [7:0] wire31 = wire28[7:0];
wire [7:0] wire32 = wire28[15:8];
wire [7:0] wire33 = wire32[7:0];
wire [3:0] wire34 = wire31[3:0];
wire [3:0] wire35 = wire31[7:4];
wire [3:0] wire36 = wire35[3:0];
wire [3:0] wire37 = wire33[3:0];
wire [3:0] wire38 = wire33[7:4];
wire [3:0] wire39 = wire38[3:0];
wire [7:0] wire40 = wire30[7:0];
wire [7:0] wire41 = wire30[15:8];
wire [7:0] wire42 = wire41[7:0];
wire [3:0] wire43 = wire40[3:0];
wire [3:0] wire44 = wire40[7:4];
wire [3:0] wire45 = wire44[3:0];
wire [3:0] wire46 = wire42[3:0];
wire [3:0] wire47 = wire42[7:4];
wire [3:0] wire48 = wire47[3:0];
wire [7:0] wire49 = {wire13, wire15};
wire [3:0] wire50 = wire49[7:4];
wire  wire51 = wire13 < wire15;
wire  wire52 = wire13 == wire15;
wire  wire53 = wire51 | wire52;
wire [3:0] wire54 = wire53 ? wire13 : wire15;
wire [3:0] wire55 = wire53 ? wire15 : wire13;
wire [7:0] wire56 = {wire54, wire55};
wire [3:0] wire57 = wire56[7:4];
wire [7:0] wire58 = {wire16, wire18};
wire [3:0] wire59 = wire58[7:4];
wire  wire60 = wire16 < wire18;
wire  wire61 = wire16 == wire18;
wire  wire62 = wire60 | wire61;
wire [3:0] wire63 = wire62 ? wire16 : wire18;
wire [3:0] wire64 = wire62 ? wire18 : wire16;
wire [7:0] wire65 = {wire63, wire64};
wire [3:0] wire66 = wire65[7:4];
wire [7:0] wire67 = {wire64, wire63};
wire [15:0] wire68 = {wire56, wire67};
wire [7:0] wire69 = wire68[15:8];
wire [3:0] wire70 = wire67[7:4];
wire  wire71 = wire54 < wire64;
wire  wire72 = wire54 == wire64;
wire  wire73 = wire71 | wire72;
wire [3:0] wire74 = wire73 ? wire54 : wire64;
wire [3:0] wire75 = wire73 ? wire64 : wire54;
wire [7:0] wire76 = {wire74, wire75};
wire [3:0] wire77 = wire76[7:4];
wire  wire78 = wire55 < wire63;
wire  wire79 = wire55 == wire63;
wire  wire80 = wire78 | wire79;
wire [3:0] wire81 = wire80 ? wire55 : wire63;
wire [3:0] wire82 = wire80 ? wire63 : wire55;
wire [7:0] wire83 = {wire81, wire82};
wire [3:0] wire84 = wire83[7:4];
wire [7:0] wire85 = {wire74, wire81};
wire [7:0] wire86 = {wire75, wire82};
wire [15:0] wire87 = {wire85, wire86};
wire [7:0] wire88 = wire87[15:8];
wire [3:0] wire89 = wire85[7:4];
wire  wire90 = wire74 < wire81;
wire  wire91 = wire74 == wire81;
wire  wire92 = wire90 | wire91;
wire [3:0] wire93 = wire92 ? wire74 : wire81;
wire [3:0] wire94 = wire92 ? wire81 : wire74;
wire [7:0] wire95 = {wire93, wire94};
wire [3:0] wire96 = wire95[7:4];
wire  wire97 = wire75 < wire82;
wire  wire98 = wire75 == wire82;
wire  wire99 = wire97 | wire98;
wire [3:0] wire100 = wire99 ? wire75 : wire82;
wire [3:0] wire101 = wire99 ? wire82 : wire75;
wire [7:0] wire102 = {wire100, wire101};
wire [3:0] wire103 = wire102[7:4];
wire [15:0] wire104 = {wire95, wire102};
wire [7:0] wire105 = {wire22, wire24};
wire [3:0] wire106 = wire105[7:4];
wire  wire107 = wire22 < wire24;
wire  wire108 = wire22 == wire24;
wire  wire109 = wire107 | wire108;
wire [3:0] wire110 = wire109 ? wire22 : wire24;
wire [3:0] wire111 = wire109 ? wire24 : wire22;
wire [7:0] wire112 = {wire110, wire111};
wire [3:0] wire113 = wire112[7:4];
wire [7:0] wire114 = {wire25, wire27};
wire [3:0] wire115 = wire114[7:4];
wire  wire116 = wire25 < wire27;
wire  wire117 = wire25 == wire27;
wire  wire118 = wire116 | wire117;
wire [3:0] wire119 = wire118 ? wire25 : wire27;
wire [3:0] wire120 = wire118 ? wire27 : wire25;
wire [7:0] wire121 = {wire119, wire120};
wire [3:0] wire122 = wire121[7:4];
wire [7:0] wire123 = {wire120, wire119};
wire [15:0] wire124 = {wire112, wire123};
wire [7:0] wire125 = wire124[15:8];
wire [3:0] wire126 = wire123[7:4];
wire  wire127 = wire110 < wire120;
wire  wire128 = wire110 == wire120;
wire  wire129 = wire127 | wire128;
wire [3:0] wire130 = wire129 ? wire110 : wire120;
wire [3:0] wire131 = wire129 ? wire120 : wire110;
wire [7:0] wire132 = {wire130, wire131};
wire [3:0] wire133 = wire132[7:4];
wire  wire134 = wire111 < wire119;
wire  wire135 = wire111 == wire119;
wire  wire136 = wire134 | wire135;
wire [3:0] wire137 = wire136 ? wire111 : wire119;
wire [3:0] wire138 = wire136 ? wire119 : wire111;
wire [7:0] wire139 = {wire137, wire138};
wire [3:0] wire140 = wire139[7:4];
wire [7:0] wire141 = {wire130, wire137};
wire [7:0] wire142 = {wire131, wire138};
wire [15:0] wire143 = {wire141, wire142};
wire [7:0] wire144 = wire143[15:8];
wire [3:0] wire145 = wire141[7:4];
wire  wire146 = wire130 < wire137;
wire  wire147 = wire130 == wire137;
wire  wire148 = wire146 | wire147;
wire [3:0] wire149 = wire148 ? wire130 : wire137;
wire [3:0] wire150 = wire148 ? wire137 : wire130;
wire [7:0] wire151 = {wire149, wire150};
wire [3:0] wire152 = wire151[7:4];
wire  wire153 = wire131 < wire138;
wire  wire154 = wire131 == wire138;
wire  wire155 = wire153 | wire154;
wire [3:0] wire156 = wire155 ? wire131 : wire138;
wire [3:0] wire157 = wire155 ? wire138 : wire131;
wire [7:0] wire158 = {wire156, wire157};
wire [3:0] wire159 = wire158[7:4];
wire [15:0] wire160 = {wire151, wire158};
wire [7:0] wire161 = wire160[15:8];
wire [7:0] wire162 = {wire157, wire156};
wire [7:0] wire163 = {wire150, wire149};
wire [15:0] wire164 = {wire162, wire163};
wire [31:0] wire165 = {wire104, wire164};
wire [15:0] wire166 = wire165[31:16];
wire [7:0] wire167 = wire104[15:8];
wire [7:0] wire168 = wire164[15:8];
wire [3:0] wire169 = wire162[7:4];
wire [3:0] wire170 = wire163[7:4];
wire  wire171 = wire93 < wire157;
wire  wire172 = wire93 == wire157;
wire  wire173 = wire171 | wire172;
wire [3:0] wire174 = wire173 ? wire93 : wire157;
wire [3:0] wire175 = wire173 ? wire157 : wire93;
wire [7:0] wire176 = {wire174, wire175};
wire [3:0] wire177 = wire176[7:4];
wire  wire178 = wire94 < wire156;
wire  wire179 = wire94 == wire156;
wire  wire180 = wire178 | wire179;
wire [3:0] wire181 = wire180 ? wire94 : wire156;
wire [3:0] wire182 = wire180 ? wire156 : wire94;
wire [7:0] wire183 = {wire181, wire182};
wire [3:0] wire184 = wire183[7:4];
wire [7:0] wire185 = {wire174, wire181};
wire [7:0] wire186 = {wire175, wire182};
wire [15:0] wire187 = {wire185, wire186};
wire [7:0] wire188 = wire187[15:8];
wire  wire189 = wire100 < wire150;
wire  wire190 = wire100 == wire150;
wire  wire191 = wire189 | wire190;
wire [3:0] wire192 = wire191 ? wire100 : wire150;
wire [3:0] wire193 = wire191 ? wire150 : wire100;
wire [7:0] wire194 = {wire192, wire193};
wire [3:0] wire195 = wire194[7:4];
wire  wire196 = wire101 < wire149;
wire  wire197 = wire101 == wire149;
wire  wire198 = wire196 | wire197;
wire [3:0] wire199 = wire198 ? wire101 : wire149;
wire [3:0] wire200 = wire198 ? wire149 : wire101;
wire [7:0] wire201 = {wire199, wire200};
wire [3:0] wire202 = wire201[7:4];
wire [7:0] wire203 = {wire192, wire199};
wire [7:0] wire204 = {wire193, wire200};
wire [15:0] wire205 = {wire203, wire204};
wire [7:0] wire206 = wire205[15:8];
wire [15:0] wire207 = {wire185, wire203};
wire [15:0] wire208 = {wire186, wire204};
wire [31:0] wire209 = {wire207, wire208};
wire [15:0] wire210 = wire209[31:16];
wire [7:0] wire211 = wire207[15:8];
wire [3:0] wire212 = wire185[7:4];
wire [3:0] wire213 = wire203[7:4];
wire  wire214 = wire174 < wire192;
wire  wire215 = wire174 == wire192;
wire  wire216 = wire214 | wire215;
wire [3:0] wire217 = wire216 ? wire174 : wire192;
wire [3:0] wire218 = wire216 ? wire192 : wire174;
wire [7:0] wire219 = {wire217, wire218};
wire [3:0] wire220 = wire219[7:4];
wire  wire221 = wire181 < wire199;
wire  wire222 = wire181 == wire199;
wire  wire223 = wire221 | wire222;
wire [3:0] wire224 = wire223 ? wire181 : wire199;
wire [3:0] wire225 = wire223 ? wire199 : wire181;
wire [7:0] wire226 = {wire224, wire225};
wire [3:0] wire227 = wire226[7:4];
wire [7:0] wire228 = {wire217, wire224};
wire [7:0] wire229 = {wire218, wire225};
wire [15:0] wire230 = {wire228, wire229};
wire [7:0] wire231 = wire230[15:8];
wire [3:0] wire232 = wire228[7:4];
wire  wire233 = wire217 < wire224;
wire  wire234 = wire217 == wire224;
wire  wire235 = wire233 | wire234;
wire [3:0] wire236 = wire235 ? wire217 : wire224;
wire [3:0] wire237 = wire235 ? wire224 : wire217;
wire [7:0] wire238 = {wire236, wire237};
wire [3:0] wire239 = wire238[7:4];
wire  wire240 = wire218 < wire225;
wire  wire241 = wire218 == wire225;
wire  wire242 = wire240 | wire241;
wire [3:0] wire243 = wire242 ? wire218 : wire225;
wire [3:0] wire244 = wire242 ? wire225 : wire218;
wire [7:0] wire245 = {wire243, wire244};
wire [3:0] wire246 = wire245[7:4];
wire [15:0] wire247 = {wire238, wire245};
wire  wire248 = wire175 < wire193;
wire  wire249 = wire175 == wire193;
wire  wire250 = wire248 | wire249;
wire [3:0] wire251 = wire250 ? wire175 : wire193;
wire [3:0] wire252 = wire250 ? wire193 : wire175;
wire [7:0] wire253 = {wire251, wire252};
wire [3:0] wire254 = wire253[7:4];
wire  wire255 = wire182 < wire200;
wire  wire256 = wire182 == wire200;
wire  wire257 = wire255 | wire256;
wire [3:0] wire258 = wire257 ? wire182 : wire200;
wire [3:0] wire259 = wire257 ? wire200 : wire182;
wire [7:0] wire260 = {wire258, wire259};
wire [3:0] wire261 = wire260[7:4];
wire [7:0] wire262 = {wire251, wire258};
wire [7:0] wire263 = {wire252, wire259};
wire [15:0] wire264 = {wire262, wire263};
wire [7:0] wire265 = wire264[15:8];
wire [3:0] wire266 = wire262[7:4];
wire  wire267 = wire251 < wire258;
wire  wire268 = wire251 == wire258;
wire  wire269 = wire267 | wire268;
wire [3:0] wire270 = wire269 ? wire251 : wire258;
wire [3:0] wire271 = wire269 ? wire258 : wire251;
wire [7:0] wire272 = {wire270, wire271};
wire [3:0] wire273 = wire272[7:4];
wire  wire274 = wire252 < wire259;
wire  wire275 = wire252 == wire259;
wire  wire276 = wire274 | wire275;
wire [3:0] wire277 = wire276 ? wire252 : wire259;
wire [3:0] wire278 = wire276 ? wire259 : wire252;
wire [7:0] wire279 = {wire277, wire278};
wire [3:0] wire280 = wire279[7:4];
wire [15:0] wire281 = {wire272, wire279};
wire [31:0] wire282 = {wire247, wire281};
wire [7:0] wire283 = {wire34, wire36};
wire [3:0] wire284 = wire283[7:4];
wire  wire285 = wire34 < wire36;
wire  wire286 = wire34 == wire36;
wire  wire287 = wire285 | wire286;
wire [3:0] wire288 = wire287 ? wire34 : wire36;
wire [3:0] wire289 = wire287 ? wire36 : wire34;
wire [7:0] wire290 = {wire288, wire289};
wire [3:0] wire291 = wire290[7:4];
wire [7:0] wire292 = {wire37, wire39};
wire [3:0] wire293 = wire292[7:4];
wire  wire294 = wire37 < wire39;
wire  wire295 = wire37 == wire39;
wire  wire296 = wire294 | wire295;
wire [3:0] wire297 = wire296 ? wire37 : wire39;
wire [3:0] wire298 = wire296 ? wire39 : wire37;
wire [7:0] wire299 = {wire297, wire298};
wire [3:0] wire300 = wire299[7:4];
wire [7:0] wire301 = {wire298, wire297};
wire [15:0] wire302 = {wire290, wire301};
wire [7:0] wire303 = wire302[15:8];
wire [3:0] wire304 = wire301[7:4];
wire  wire305 = wire288 < wire298;
wire  wire306 = wire288 == wire298;
wire  wire307 = wire305 | wire306;
wire [3:0] wire308 = wire307 ? wire288 : wire298;
wire [3:0] wire309 = wire307 ? wire298 : wire288;
wire [7:0] wire310 = {wire308, wire309};
wire [3:0] wire311 = wire310[7:4];
wire  wire312 = wire289 < wire297;
wire  wire313 = wire289 == wire297;
wire  wire314 = wire312 | wire313;
wire [3:0] wire315 = wire314 ? wire289 : wire297;
wire [3:0] wire316 = wire314 ? wire297 : wire289;
wire [7:0] wire317 = {wire315, wire316};
wire [3:0] wire318 = wire317[7:4];
wire [7:0] wire319 = {wire308, wire315};
wire [7:0] wire320 = {wire309, wire316};
wire [15:0] wire321 = {wire319, wire320};
wire [7:0] wire322 = wire321[15:8];
wire [3:0] wire323 = wire319[7:4];
wire  wire324 = wire308 < wire315;
wire  wire325 = wire308 == wire315;
wire  wire326 = wire324 | wire325;
wire [3:0] wire327 = wire326 ? wire308 : wire315;
wire [3:0] wire328 = wire326 ? wire315 : wire308;
wire [7:0] wire329 = {wire327, wire328};
wire [3:0] wire330 = wire329[7:4];
wire  wire331 = wire309 < wire316;
wire  wire332 = wire309 == wire316;
wire  wire333 = wire331 | wire332;
wire [3:0] wire334 = wire333 ? wire309 : wire316;
wire [3:0] wire335 = wire333 ? wire316 : wire309;
wire [7:0] wire336 = {wire334, wire335};
wire [3:0] wire337 = wire336[7:4];
wire [15:0] wire338 = {wire329, wire336};
wire [7:0] wire339 = {wire43, wire45};
wire [3:0] wire340 = wire339[7:4];
wire  wire341 = wire43 < wire45;
wire  wire342 = wire43 == wire45;
wire  wire343 = wire341 | wire342;
wire [3:0] wire344 = wire343 ? wire43 : wire45;
wire [3:0] wire345 = wire343 ? wire45 : wire43;
wire [7:0] wire346 = {wire344, wire345};
wire [3:0] wire347 = wire346[7:4];
wire [7:0] wire348 = {wire46, wire48};
wire [3:0] wire349 = wire348[7:4];
wire  wire350 = wire46 < wire48;
wire  wire351 = wire46 == wire48;
wire  wire352 = wire350 | wire351;
wire [3:0] wire353 = wire352 ? wire46 : wire48;
wire [3:0] wire354 = wire352 ? wire48 : wire46;
wire [7:0] wire355 = {wire353, wire354};
wire [3:0] wire356 = wire355[7:4];
wire [7:0] wire357 = {wire354, wire353};
wire [15:0] wire358 = {wire346, wire357};
wire [7:0] wire359 = wire358[15:8];
wire [3:0] wire360 = wire357[7:4];
wire  wire361 = wire344 < wire354;
wire  wire362 = wire344 == wire354;
wire  wire363 = wire361 | wire362;
wire [3:0] wire364 = wire363 ? wire344 : wire354;
wire [3:0] wire365 = wire363 ? wire354 : wire344;
wire [7:0] wire366 = {wire364, wire365};
wire [3:0] wire367 = wire366[7:4];
wire  wire368 = wire345 < wire353;
wire  wire369 = wire345 == wire353;
wire  wire370 = wire368 | wire369;
wire [3:0] wire371 = wire370 ? wire345 : wire353;
wire [3:0] wire372 = wire370 ? wire353 : wire345;
wire [7:0] wire373 = {wire371, wire372};
wire [3:0] wire374 = wire373[7:4];
wire [7:0] wire375 = {wire364, wire371};
wire [7:0] wire376 = {wire365, wire372};
wire [15:0] wire377 = {wire375, wire376};
wire [7:0] wire378 = wire377[15:8];
wire [3:0] wire379 = wire375[7:4];
wire  wire380 = wire364 < wire371;
wire  wire381 = wire364 == wire371;
wire  wire382 = wire380 | wire381;
wire [3:0] wire383 = wire382 ? wire364 : wire371;
wire [3:0] wire384 = wire382 ? wire371 : wire364;
wire [7:0] wire385 = {wire383, wire384};
wire [3:0] wire386 = wire385[7:4];
wire  wire387 = wire365 < wire372;
wire  wire388 = wire365 == wire372;
wire  wire389 = wire387 | wire388;
wire [3:0] wire390 = wire389 ? wire365 : wire372;
wire [3:0] wire391 = wire389 ? wire372 : wire365;
wire [7:0] wire392 = {wire390, wire391};
wire [3:0] wire393 = wire392[7:4];
wire [15:0] wire394 = {wire385, wire392};
wire [7:0] wire395 = wire394[15:8];
wire [7:0] wire396 = {wire391, wire390};
wire [7:0] wire397 = {wire384, wire383};
wire [15:0] wire398 = {wire396, wire397};
wire [31:0] wire399 = {wire338, wire398};
wire [15:0] wire400 = wire399[31:16];
wire [7:0] wire401 = wire338[15:8];
wire [7:0] wire402 = wire398[15:8];
wire [3:0] wire403 = wire396[7:4];
wire [3:0] wire404 = wire397[7:4];
wire  wire405 = wire327 < wire391;
wire  wire406 = wire327 == wire391;
wire  wire407 = wire405 | wire406;
wire [3:0] wire408 = wire407 ? wire327 : wire391;
wire [3:0] wire409 = wire407 ? wire391 : wire327;
wire [7:0] wire410 = {wire408, wire409};
wire [3:0] wire411 = wire410[7:4];
wire  wire412 = wire328 < wire390;
wire  wire413 = wire328 == wire390;
wire  wire414 = wire412 | wire413;
wire [3:0] wire415 = wire414 ? wire328 : wire390;
wire [3:0] wire416 = wire414 ? wire390 : wire328;
wire [7:0] wire417 = {wire415, wire416};
wire [3:0] wire418 = wire417[7:4];
wire [7:0] wire419 = {wire408, wire415};
wire [7:0] wire420 = {wire409, wire416};
wire [15:0] wire421 = {wire419, wire420};
wire [7:0] wire422 = wire421[15:8];
wire  wire423 = wire334 < wire384;
wire  wire424 = wire334 == wire384;
wire  wire425 = wire423 | wire424;
wire [3:0] wire426 = wire425 ? wire334 : wire384;
wire [3:0] wire427 = wire425 ? wire384 : wire334;
wire [7:0] wire428 = {wire426, wire427};
wire [3:0] wire429 = wire428[7:4];
wire  wire430 = wire335 < wire383;
wire  wire431 = wire335 == wire383;
wire  wire432 = wire430 | wire431;
wire [3:0] wire433 = wire432 ? wire335 : wire383;
wire [3:0] wire434 = wire432 ? wire383 : wire335;
wire [7:0] wire435 = {wire433, wire434};
wire [3:0] wire436 = wire435[7:4];
wire [7:0] wire437 = {wire426, wire433};
wire [7:0] wire438 = {wire427, wire434};
wire [15:0] wire439 = {wire437, wire438};
wire [7:0] wire440 = wire439[15:8];
wire [15:0] wire441 = {wire419, wire437};
wire [15:0] wire442 = {wire420, wire438};
wire [31:0] wire443 = {wire441, wire442};
wire [15:0] wire444 = wire443[31:16];
wire [7:0] wire445 = wire441[15:8];
wire [3:0] wire446 = wire419[7:4];
wire [3:0] wire447 = wire437[7:4];
wire  wire448 = wire408 < wire426;
wire  wire449 = wire408 == wire426;
wire  wire450 = wire448 | wire449;
wire [3:0] wire451 = wire450 ? wire408 : wire426;
wire [3:0] wire452 = wire450 ? wire426 : wire408;
wire [7:0] wire453 = {wire451, wire452};
wire [3:0] wire454 = wire453[7:4];
wire  wire455 = wire415 < wire433;
wire  wire456 = wire415 == wire433;
wire  wire457 = wire455 | wire456;
wire [3:0] wire458 = wire457 ? wire415 : wire433;
wire [3:0] wire459 = wire457 ? wire433 : wire415;
wire [7:0] wire460 = {wire458, wire459};
wire [3:0] wire461 = wire460[7:4];
wire [7:0] wire462 = {wire451, wire458};
wire [7:0] wire463 = {wire452, wire459};
wire [15:0] wire464 = {wire462, wire463};
wire [7:0] wire465 = wire464[15:8];
wire [3:0] wire466 = wire462[7:4];
wire  wire467 = wire451 < wire458;
wire  wire468 = wire451 == wire458;
wire  wire469 = wire467 | wire468;
wire [3:0] wire470 = wire469 ? wire451 : wire458;
wire [3:0] wire471 = wire469 ? wire458 : wire451;
wire [7:0] wire472 = {wire470, wire471};
wire [3:0] wire473 = wire472[7:4];
wire  wire474 = wire452 < wire459;
wire  wire475 = wire452 == wire459;
wire  wire476 = wire474 | wire475;
wire [3:0] wire477 = wire476 ? wire452 : wire459;
wire [3:0] wire478 = wire476 ? wire459 : wire452;
wire [7:0] wire479 = {wire477, wire478};
wire [3:0] wire480 = wire479[7:4];
wire [15:0] wire481 = {wire472, wire479};
wire  wire482 = wire409 < wire427;
wire  wire483 = wire409 == wire427;
wire  wire484 = wire482 | wire483;
wire [3:0] wire485 = wire484 ? wire409 : wire427;
wire [3:0] wire486 = wire484 ? wire427 : wire409;
wire [7:0] wire487 = {wire485, wire486};
wire [3:0] wire488 = wire487[7:4];
wire  wire489 = wire416 < wire434;
wire  wire490 = wire416 == wire434;
wire  wire491 = wire489 | wire490;
wire [3:0] wire492 = wire491 ? wire416 : wire434;
wire [3:0] wire493 = wire491 ? wire434 : wire416;
wire [7:0] wire494 = {wire492, wire493};
wire [3:0] wire495 = wire494[7:4];
wire [7:0] wire496 = {wire485, wire492};
wire [7:0] wire497 = {wire486, wire493};
wire [15:0] wire498 = {wire496, wire497};
wire [7:0] wire499 = wire498[15:8];
wire [3:0] wire500 = wire496[7:4];
wire  wire501 = wire485 < wire492;
wire  wire502 = wire485 == wire492;
wire  wire503 = wire501 | wire502;
wire [3:0] wire504 = wire503 ? wire485 : wire492;
wire [3:0] wire505 = wire503 ? wire492 : wire485;
wire [7:0] wire506 = {wire504, wire505};
wire [3:0] wire507 = wire506[7:4];
wire  wire508 = wire486 < wire493;
wire  wire509 = wire486 == wire493;
wire  wire510 = wire508 | wire509;
wire [3:0] wire511 = wire510 ? wire486 : wire493;
wire [3:0] wire512 = wire510 ? wire493 : wire486;
wire [7:0] wire513 = {wire511, wire512};
wire [3:0] wire514 = wire513[7:4];
wire [15:0] wire515 = {wire506, wire513};
wire [31:0] wire516 = {wire481, wire515};
wire [15:0] wire517 = wire516[31:16];
wire [7:0] wire518 = wire481[15:8];
wire [7:0] wire519 = wire515[15:8];
wire [7:0] wire520 = {wire512, wire511};
wire [7:0] wire521 = {wire505, wire504};
wire [15:0] wire522 = {wire520, wire521};
wire [7:0] wire523 = {wire478, wire477};
wire [7:0] wire524 = {wire471, wire470};
wire [15:0] wire525 = {wire523, wire524};
wire [31:0] wire526 = {wire522, wire525};
wire [63:0] wire527 = {wire282, wire526};
wire [31:0] wire528 = wire527[63:32];
wire [15:0] wire529 = wire282[31:16];
wire [7:0] wire530 = wire247[15:8];
wire [7:0] wire531 = wire281[15:8];
wire [15:0] wire532 = wire526[31:16];
wire [7:0] wire533 = wire522[15:8];
wire [3:0] wire534 = wire520[7:4];
wire [3:0] wire535 = wire521[7:4];
wire [7:0] wire536 = wire525[15:8];
wire [3:0] wire537 = wire523[7:4];
wire [3:0] wire538 = wire524[7:4];
wire  wire539 = wire236 < wire512;
wire  wire540 = wire236 == wire512;
wire  wire541 = wire539 | wire540;
wire [3:0] wire542 = wire541 ? wire236 : wire512;
wire [3:0] wire543 = wire541 ? wire512 : wire236;
wire [7:0] wire544 = {wire542, wire543};
wire [3:0] wire545 = wire544[7:4];
wire  wire546 = wire237 < wire511;
wire  wire547 = wire237 == wire511;
wire  wire548 = wire546 | wire547;
wire [3:0] wire549 = wire548 ? wire237 : wire511;
wire [3:0] wire550 = wire548 ? wire511 : wire237;
wire [7:0] wire551 = {wire549, wire550};
wire [3:0] wire552 = wire551[7:4];
wire [7:0] wire553 = {wire542, wire549};
wire [7:0] wire554 = {wire543, wire550};
wire [15:0] wire555 = {wire553, wire554};
wire [7:0] wire556 = wire555[15:8];
wire  wire557 = wire243 < wire505;
wire  wire558 = wire243 == wire505;
wire  wire559 = wire557 | wire558;
wire [3:0] wire560 = wire559 ? wire243 : wire505;
wire [3:0] wire561 = wire559 ? wire505 : wire243;
wire [7:0] wire562 = {wire560, wire561};
wire [3:0] wire563 = wire562[7:4];
wire  wire564 = wire244 < wire504;
wire  wire565 = wire244 == wire504;
wire  wire566 = wire564 | wire565;
wire [3:0] wire567 = wire566 ? wire244 : wire504;
wire [3:0] wire568 = wire566 ? wire504 : wire244;
wire [7:0] wire569 = {wire567, wire568};
wire [3:0] wire570 = wire569[7:4];
wire [7:0] wire571 = {wire560, wire567};
wire [7:0] wire572 = {wire561, wire568};
wire [15:0] wire573 = {wire571, wire572};
wire [7:0] wire574 = wire573[15:8];
wire [15:0] wire575 = {wire553, wire571};
wire [15:0] wire576 = {wire554, wire572};
wire [31:0] wire577 = {wire575, wire576};
wire [15:0] wire578 = wire577[31:16];
wire  wire579 = wire270 < wire478;
wire  wire580 = wire270 == wire478;
wire  wire581 = wire579 | wire580;
wire [3:0] wire582 = wire581 ? wire270 : wire478;
wire [3:0] wire583 = wire581 ? wire478 : wire270;
wire [7:0] wire584 = {wire582, wire583};
wire [3:0] wire585 = wire584[7:4];
wire  wire586 = wire271 < wire477;
wire  wire587 = wire271 == wire477;
wire  wire588 = wire586 | wire587;
wire [3:0] wire589 = wire588 ? wire271 : wire477;
wire [3:0] wire590 = wire588 ? wire477 : wire271;
wire [7:0] wire591 = {wire589, wire590};
wire [3:0] wire592 = wire591[7:4];
wire [7:0] wire593 = {wire582, wire589};
wire [7:0] wire594 = {wire583, wire590};
wire [15:0] wire595 = {wire593, wire594};
wire [7:0] wire596 = wire595[15:8];
wire  wire597 = wire277 < wire471;
wire  wire598 = wire277 == wire471;
wire  wire599 = wire597 | wire598;
wire [3:0] wire600 = wire599 ? wire277 : wire471;
wire [3:0] wire601 = wire599 ? wire471 : wire277;
wire [7:0] wire602 = {wire600, wire601};
wire [3:0] wire603 = wire602[7:4];
wire  wire604 = wire278 < wire470;
wire  wire605 = wire278 == wire470;
wire  wire606 = wire604 | wire605;
wire [3:0] wire607 = wire606 ? wire278 : wire470;
wire [3:0] wire608 = wire606 ? wire470 : wire278;
wire [7:0] wire609 = {wire607, wire608};
wire [3:0] wire610 = wire609[7:4];
wire [7:0] wire611 = {wire600, wire607};
wire [7:0] wire612 = {wire601, wire608};
wire [15:0] wire613 = {wire611, wire612};
wire [7:0] wire614 = wire613[15:8];
wire [15:0] wire615 = {wire593, wire611};
wire [15:0] wire616 = {wire594, wire612};
wire [31:0] wire617 = {wire615, wire616};
wire [15:0] wire618 = wire617[31:16];
wire [31:0] wire619 = {wire575, wire615};
wire [31:0] wire620 = {wire576, wire616};
wire [63:0] wire621 = {wire619, wire620};
wire [31:0] wire622 = wire621[63:32];
wire [15:0] wire623 = wire619[31:16];
wire [7:0] wire624 = wire575[15:8];
wire [3:0] wire625 = wire553[7:4];
wire [3:0] wire626 = wire571[7:4];
wire [7:0] wire627 = wire615[15:8];
wire [3:0] wire628 = wire593[7:4];
wire [3:0] wire629 = wire611[7:4];
wire  wire630 = wire542 < wire582;
wire  wire631 = wire542 == wire582;
wire  wire632 = wire630 | wire631;
wire [3:0] wire633 = wire632 ? wire542 : wire582;
wire [3:0] wire634 = wire632 ? wire582 : wire542;
wire [7:0] wire635 = {wire633, wire634};
wire [3:0] wire636 = wire635[7:4];
wire  wire637 = wire549 < wire589;
wire  wire638 = wire549 == wire589;
wire  wire639 = wire637 | wire638;
wire [3:0] wire640 = wire639 ? wire549 : wire589;
wire [3:0] wire641 = wire639 ? wire589 : wire549;
wire [7:0] wire642 = {wire640, wire641};
wire [3:0] wire643 = wire642[7:4];
wire [7:0] wire644 = {wire633, wire640};
wire [7:0] wire645 = {wire634, wire641};
wire [15:0] wire646 = {wire644, wire645};
wire [7:0] wire647 = wire646[15:8];
wire  wire648 = wire560 < wire600;
wire  wire649 = wire560 == wire600;
wire  wire650 = wire648 | wire649;
wire [3:0] wire651 = wire650 ? wire560 : wire600;
wire [3:0] wire652 = wire650 ? wire600 : wire560;
wire [7:0] wire653 = {wire651, wire652};
wire [3:0] wire654 = wire653[7:4];
wire  wire655 = wire567 < wire607;
wire  wire656 = wire567 == wire607;
wire  wire657 = wire655 | wire656;
wire [3:0] wire658 = wire657 ? wire567 : wire607;
wire [3:0] wire659 = wire657 ? wire607 : wire567;
wire [7:0] wire660 = {wire658, wire659};
wire [3:0] wire661 = wire660[7:4];
wire [7:0] wire662 = {wire651, wire658};
wire [7:0] wire663 = {wire652, wire659};
wire [15:0] wire664 = {wire662, wire663};
wire [7:0] wire665 = wire664[15:8];
wire [15:0] wire666 = {wire644, wire662};
wire [15:0] wire667 = {wire645, wire663};
wire [31:0] wire668 = {wire666, wire667};
wire [15:0] wire669 = wire668[31:16];
wire [7:0] wire670 = wire666[15:8];
wire [3:0] wire671 = wire644[7:4];
wire [3:0] wire672 = wire662[7:4];
wire  wire673 = wire633 < wire651;
wire  wire674 = wire633 == wire651;
wire  wire675 = wire673 | wire674;
wire [3:0] wire676 = wire675 ? wire633 : wire651;
wire [3:0] wire677 = wire675 ? wire651 : wire633;
wire [7:0] wire678 = {wire676, wire677};
wire [3:0] wire679 = wire678[7:4];
wire  wire680 = wire640 < wire658;
wire  wire681 = wire640 == wire658;
wire  wire682 = wire680 | wire681;
wire [3:0] wire683 = wire682 ? wire640 : wire658;
wire [3:0] wire684 = wire682 ? wire658 : wire640;
wire [7:0] wire685 = {wire683, wire684};
wire [3:0] wire686 = wire685[7:4];
wire [7:0] wire687 = {wire676, wire683};
wire [7:0] wire688 = {wire677, wire684};
wire [15:0] wire689 = {wire687, wire688};
wire [7:0] wire690 = wire689[15:8];
wire [3:0] wire691 = wire687[7:4];
wire  wire692 = wire676 < wire683;
wire  wire693 = wire676 == wire683;
wire  wire694 = wire692 | wire693;
wire [3:0] wire695 = wire694 ? wire676 : wire683;
wire [3:0] wire696 = wire694 ? wire683 : wire676;
wire [7:0] wire697 = {wire695, wire696};
wire [3:0] wire698 = wire697[7:4];
wire  wire699 = wire677 < wire684;
wire  wire700 = wire677 == wire684;
wire  wire701 = wire699 | wire700;
wire [3:0] wire702 = wire701 ? wire677 : wire684;
wire [3:0] wire703 = wire701 ? wire684 : wire677;
wire [7:0] wire704 = {wire702, wire703};
wire [3:0] wire705 = wire704[7:4];
wire [15:0] wire706 = {wire697, wire704};
wire  wire707 = wire634 < wire652;
wire  wire708 = wire634 == wire652;
wire  wire709 = wire707 | wire708;
wire [3:0] wire710 = wire709 ? wire634 : wire652;
wire [3:0] wire711 = wire709 ? wire652 : wire634;
wire [7:0] wire712 = {wire710, wire711};
wire [3:0] wire713 = wire712[7:4];
wire  wire714 = wire641 < wire659;
wire  wire715 = wire641 == wire659;
wire  wire716 = wire714 | wire715;
wire [3:0] wire717 = wire716 ? wire641 : wire659;
wire [3:0] wire718 = wire716 ? wire659 : wire641;
wire [7:0] wire719 = {wire717, wire718};
wire [3:0] wire720 = wire719[7:4];
wire [7:0] wire721 = {wire710, wire717};
wire [7:0] wire722 = {wire711, wire718};
wire [15:0] wire723 = {wire721, wire722};
wire [7:0] wire724 = wire723[15:8];
wire [3:0] wire725 = wire721[7:4];
wire  wire726 = wire710 < wire717;
wire  wire727 = wire710 == wire717;
wire  wire728 = wire726 | wire727;
wire [3:0] wire729 = wire728 ? wire710 : wire717;
wire [3:0] wire730 = wire728 ? wire717 : wire710;
wire [7:0] wire731 = {wire729, wire730};
wire [3:0] wire732 = wire731[7:4];
wire  wire733 = wire711 < wire718;
wire  wire734 = wire711 == wire718;
wire  wire735 = wire733 | wire734;
wire [3:0] wire736 = wire735 ? wire711 : wire718;
wire [3:0] wire737 = wire735 ? wire718 : wire711;
wire [7:0] wire738 = {wire736, wire737};
wire [3:0] wire739 = wire738[7:4];
wire [15:0] wire740 = {wire731, wire738};
wire [31:0] wire741 = {wire706, wire740};
wire  wire742 = wire543 < wire583;
wire  wire743 = wire543 == wire583;
wire  wire744 = wire742 | wire743;
wire [3:0] wire745 = wire744 ? wire543 : wire583;
wire [3:0] wire746 = wire744 ? wire583 : wire543;
wire [7:0] wire747 = {wire745, wire746};
wire [3:0] wire748 = wire747[7:4];
wire  wire749 = wire550 < wire590;
wire  wire750 = wire550 == wire590;
wire  wire751 = wire749 | wire750;
wire [3:0] wire752 = wire751 ? wire550 : wire590;
wire [3:0] wire753 = wire751 ? wire590 : wire550;
wire [7:0] wire754 = {wire752, wire753};
wire [3:0] wire755 = wire754[7:4];
wire [7:0] wire756 = {wire745, wire752};
wire [7:0] wire757 = {wire746, wire753};
wire [15:0] wire758 = {wire756, wire757};
wire [7:0] wire759 = wire758[15:8];
wire  wire760 = wire561 < wire601;
wire  wire761 = wire561 == wire601;
wire  wire762 = wire760 | wire761;
wire [3:0] wire763 = wire762 ? wire561 : wire601;
wire [3:0] wire764 = wire762 ? wire601 : wire561;
wire [7:0] wire765 = {wire763, wire764};
wire [3:0] wire766 = wire765[7:4];
wire  wire767 = wire568 < wire608;
wire  wire768 = wire568 == wire608;
wire  wire769 = wire767 | wire768;
wire [3:0] wire770 = wire769 ? wire568 : wire608;
wire [3:0] wire771 = wire769 ? wire608 : wire568;
wire [7:0] wire772 = {wire770, wire771};
wire [3:0] wire773 = wire772[7:4];
wire [7:0] wire774 = {wire763, wire770};
wire [7:0] wire775 = {wire764, wire771};
wire [15:0] wire776 = {wire774, wire775};
wire [7:0] wire777 = wire776[15:8];
wire [15:0] wire778 = {wire756, wire774};
wire [15:0] wire779 = {wire757, wire775};
wire [31:0] wire780 = {wire778, wire779};
wire [15:0] wire781 = wire780[31:16];
wire [7:0] wire782 = wire778[15:8];
wire [3:0] wire783 = wire756[7:4];
wire [3:0] wire784 = wire774[7:4];
wire  wire785 = wire745 < wire763;
wire  wire786 = wire745 == wire763;
wire  wire787 = wire785 | wire786;
wire [3:0] wire788 = wire787 ? wire745 : wire763;
wire [3:0] wire789 = wire787 ? wire763 : wire745;
wire [7:0] wire790 = {wire788, wire789};
wire [3:0] wire791 = wire790[7:4];
wire  wire792 = wire752 < wire770;
wire  wire793 = wire752 == wire770;
wire  wire794 = wire792 | wire793;
wire [3:0] wire795 = wire794 ? wire752 : wire770;
wire [3:0] wire796 = wire794 ? wire770 : wire752;
wire [7:0] wire797 = {wire795, wire796};
wire [3:0] wire798 = wire797[7:4];
wire [7:0] wire799 = {wire788, wire795};
wire [7:0] wire800 = {wire789, wire796};
wire [15:0] wire801 = {wire799, wire800};
wire [7:0] wire802 = wire801[15:8];
wire [3:0] wire803 = wire799[7:4];
wire  wire804 = wire788 < wire795;
wire  wire805 = wire788 == wire795;
wire  wire806 = wire804 | wire805;
wire [3:0] wire807 = wire806 ? wire788 : wire795;
wire [3:0] wire808 = wire806 ? wire795 : wire788;
wire [7:0] wire809 = {wire807, wire808};
wire [3:0] wire810 = wire809[7:4];
wire  wire811 = wire789 < wire796;
wire  wire812 = wire789 == wire796;
wire  wire813 = wire811 | wire812;
wire [3:0] wire814 = wire813 ? wire789 : wire796;
wire [3:0] wire815 = wire813 ? wire796 : wire789;
wire [7:0] wire816 = {wire814, wire815};
wire [3:0] wire817 = wire816[7:4];
wire [15:0] wire818 = {wire809, wire816};
wire  wire819 = wire746 < wire764;
wire  wire820 = wire746 == wire764;
wire  wire821 = wire819 | wire820;
wire [3:0] wire822 = wire821 ? wire746 : wire764;
wire [3:0] wire823 = wire821 ? wire764 : wire746;
wire [7:0] wire824 = {wire822, wire823};
wire [3:0] wire825 = wire824[7:4];
wire  wire826 = wire753 < wire771;
wire  wire827 = wire753 == wire771;
wire  wire828 = wire826 | wire827;
wire [3:0] wire829 = wire828 ? wire753 : wire771;
wire [3:0] wire830 = wire828 ? wire771 : wire753;
wire [7:0] wire831 = {wire829, wire830};
wire [3:0] wire832 = wire831[7:4];
wire [7:0] wire833 = {wire822, wire829};
wire [7:0] wire834 = {wire823, wire830};
wire [15:0] wire835 = {wire833, wire834};
wire [7:0] wire836 = wire835[15:8];
wire [3:0] wire837 = wire833[7:4];
wire  wire838 = wire822 < wire829;
wire  wire839 = wire822 == wire829;
wire  wire840 = wire838 | wire839;
wire [3:0] wire841 = wire840 ? wire822 : wire829;
wire [3:0] wire842 = wire840 ? wire829 : wire822;
wire [7:0] wire843 = {wire841, wire842};
wire [3:0] wire844 = wire843[7:4];
wire  wire845 = wire823 < wire830;
wire  wire846 = wire823 == wire830;
wire  wire847 = wire845 | wire846;
wire [3:0] wire848 = wire847 ? wire823 : wire830;
wire [3:0] wire849 = wire847 ? wire830 : wire823;
wire [7:0] wire850 = {wire848, wire849};
wire [3:0] wire851 = wire850[7:4];
wire [15:0] wire852 = {wire843, wire850};
wire [31:0] wire853 = {wire818, wire852};
wire [63:0] wire854 = {wire741, wire853};
// effects 
assign guard = wire1;
assign value = wire854;
always@(posedge clk)
begin
	if(rst_n)
		begin
// reset 
		end
	else
		begin
	if(wire1)
		begin
// put  debug code here (display, stop, ...)
		end
		end
end
endmodule
