module Stack (clk, rst_n, guard, value);
integer index; // Used for initialisations
input clk;
input rst_n;
output guard;
output [-1:0] value;
// state declarations
reg [11:0] reg_0 [255:0];
reg [7:0] reg_1;
reg [7:0] reg_2 [255:0];
reg [7:0] reg_3;
reg [7:0] reg_4 [255:0];
// bindings 
wire  wire0 = 0'b0;
wire  wire1 = 1'b1;
wire  wire2 = 1'b0;
wire [7:0] wire3 = reg_1;
wire [11:0] wire4 = reg_0[wire3];
wire [3:0] wire5 = wire4[3:0];
wire [3:0] wire6 = 4'b0;
wire  wire7 = wire5 == wire6;
wire [7:0] wire8 = reg_3;
wire [7:0] wire9 = wire4[11:4];
wire [7:0] wire10 = 8'b1;
wire [7:0] wire11 = wire8 + wire10;
wire [7:0] wire12 = wire3 + wire10;
wire [3:0] wire13 = wire4[3:0];
wire  wire14 = wire13 == wire6;
wire  wire15 = ~ wire14;
wire [3:0] wire16 = wire4[3:0];
wire [3:0] wire17 = 4'b1;
wire  wire18 = wire16 == wire17;
wire [7:0] wire19 = wire4[11:4];
wire [7:0] wire20 = reg_4[wire19];
wire [3:0] wire21 = wire4[3:0];
wire  wire22 = wire21 == wire17;
wire  wire23 = ~ wire22;
wire [3:0] wire24 = wire4[3:0];
wire [3:0] wire25 = 4'b10;
wire  wire26 = wire24 == wire25;
wire [7:0] wire27 = wire8 - wire10;
wire [7:0] wire28 = reg_2[wire27];
wire [7:0] wire29 = wire4[11:4];
wire [3:0] wire30 = wire4[3:0];
wire  wire31 = wire30 == wire25;
wire  wire32 = ~ wire31;
wire [3:0] wire33 = wire4[3:0];
wire [3:0] wire34 = 4'b11;
wire  wire35 = wire33 == wire34;
wire [7:0] wire36 = reg_2[wire27];
wire [7:0] wire37 = 8'b10;
wire [7:0] wire38 = wire8 - wire37;
wire [7:0] wire39 = reg_2[wire38];
wire [7:0] wire40 = wire39 + wire36;
wire [3:0] wire41 = wire4[3:0];
wire  wire42 = wire41 == wire34;
wire  wire43 = ~ wire42;
wire [3:0] wire44 = wire4[3:0];
wire [3:0] wire45 = 4'b100;
wire  wire46 = wire44 == wire45;
wire [7:0] wire47 = reg_2[wire27];
wire [7:0] wire48 = reg_2[wire38];
wire [7:0] wire49 = wire48 - wire47;
wire [3:0] wire50 = wire4[3:0];
wire  wire51 = wire50 == wire45;
wire  wire52 = ~ wire51;
wire [3:0] wire53 = wire4[3:0];
wire [3:0] wire54 = 4'b101;
wire  wire55 = wire53 == wire54;
wire [7:0] wire56 = wire4[11:4];
wire [7:0] wire57 = wire12 + wire56;
wire [3:0] wire58 = wire4[3:0];
wire  wire59 = wire58 == wire54;
wire  wire60 = ~ wire59;
wire [3:0] wire61 = wire4[3:0];
wire [3:0] wire62 = 4'b110;
wire  wire63 = wire61 == wire62;
wire [7:0] wire64 = wire4[11:4];
wire [7:0] wire65 = wire12 - wire64;
wire [3:0] wire66 = wire4[3:0];
wire  wire67 = wire66 == wire62;
wire  wire68 = ~ wire67;
wire [3:0] wire69 = wire4[3:0];
wire [3:0] wire70 = 4'b111;
wire  wire71 = wire69 == wire70;
wire [7:0] wire72 = reg_2[wire27];
wire [7:0] wire73 = reg_2[wire38];
wire  wire74 = wire73 == wire72;
wire [7:0] wire75 = wire4[11:4];
wire [7:0] wire76 = wire12 + wire75;
wire [3:0] wire77 = wire4[3:0];
wire  wire78 = wire77 == wire70;
wire  wire79 = ~ wire78;
wire [3:0] wire80 = wire4[3:0];
wire [3:0] wire81 = 4'b1000;
wire  wire82 = wire80 == wire81;
wire [7:0] wire83 = reg_2[wire27];
wire [7:0] wire84 = reg_2[wire38];
wire  wire85 = wire84 == wire83;
wire  wire86 = ~ wire85;
wire [7:0] wire87 = wire4[11:4];
wire [7:0] wire88 = wire12 + wire87;
wire [3:0] wire89 = wire4[3:0];
wire  wire90 = wire89 == wire81;
wire  wire91 = ~ wire90;
wire [3:0] wire92 = wire4[3:0];
wire [3:0] wire93 = 4'b1001;
wire  wire94 = wire92 == wire93;
wire [7:0] wire95 = reg_2[wire27];
wire [7:0] wire96 = reg_2[wire38];
wire  wire97 = wire96 < wire95;
wire  wire98 = wire96 == wire95;
wire  wire99 = wire97 | wire98;
wire [7:0] wire100 = wire4[11:4];
wire [7:0] wire101 = wire12 + wire100;
wire [3:0] wire102 = wire4[3:0];
wire  wire103 = wire102 == wire93;
wire  wire104 = ~ wire103;
wire [3:0] wire105 = wire4[3:0];
wire [3:0] wire106 = 4'b1010;
wire  wire107 = wire105 == wire106;
wire [7:0] wire108 = reg_2[wire27];
wire [7:0] wire109 = reg_2[wire38];
wire  wire110 = wire108 < wire109;
wire [7:0] wire111 = wire4[11:4];
wire [7:0] wire112 = wire12 + wire111;
wire [3:0] wire113 = wire4[3:0];
wire  wire114 = wire113 == wire106;
wire  wire115 = ~ wire114;
wire  wire116 = wire107 | wire115;
wire  wire117 = wire104 & wire116;
wire  wire118 = wire94 | wire117;
wire  wire119 = wire91 & wire118;
wire  wire120 = wire82 | wire119;
wire  wire121 = wire79 & wire120;
wire  wire122 = wire71 | wire121;
wire  wire123 = wire68 & wire122;
wire  wire124 = wire63 | wire123;
wire  wire125 = wire60 & wire124;
wire  wire126 = wire55 | wire125;
wire  wire127 = wire52 & wire126;
wire  wire128 = wire46 | wire127;
wire  wire129 = wire43 & wire128;
wire  wire130 = wire35 | wire129;
wire  wire131 = wire32 & wire130;
wire  wire132 = wire26 | wire131;
wire  wire133 = wire23 & wire132;
wire  wire134 = wire18 | wire133;
wire  wire135 = wire15 & wire134;
wire  wire136 = wire7 | wire135;
wire  wire137 = wire136 & wire7;
wire  wire138 = ~ wire7;
wire  wire139 = wire138 & wire135;
wire  wire140 = wire139 & wire18;
wire  wire141 = wire137 | wire140;
wire [7:0] wire142 = wire137 ? wire9 : wire20;
wire  wire143 = ~ wire18;
wire  wire144 = wire143 & wire133;
wire  wire145 = wire139 & wire144;
wire  wire146 = wire145 & wire26;
wire  wire147 = wire141 | wire146;
wire [7:0] wire148 = wire141 ? wire11 : wire27;
wire  wire149 = ~ wire26;
wire  wire150 = wire149 & wire131;
wire  wire151 = wire145 & wire150;
wire  wire152 = wire151 & wire35;
wire  wire153 = wire141 | wire152;
wire [7:0] wire154 = wire141 ? wire8 : wire38;
wire [7:0] wire155 = wire141 ? wire142 : wire40;
wire  wire156 = wire147 | wire152;
wire [7:0] wire157 = wire147 ? wire148 : wire27;
wire  wire158 = ~ wire35;
wire  wire159 = wire158 & wire129;
wire  wire160 = wire151 & wire159;
wire  wire161 = wire160 & wire46;
wire  wire162 = wire153 | wire161;
wire [7:0] wire163 = wire153 ? wire154 : wire38;
wire [7:0] wire164 = wire153 ? wire155 : wire49;
wire  wire165 = wire156 | wire161;
wire [7:0] wire166 = wire156 ? wire157 : wire27;
wire  wire167 = ~ wire46;
wire  wire168 = wire167 & wire127;
wire  wire169 = wire160 & wire168;
wire  wire170 = wire169 & wire55;
wire  wire171 = wire165 | wire170;
wire [7:0] wire172 = wire165 ? wire12 : wire57;
wire  wire173 = ~ wire55;
wire  wire174 = wire173 & wire125;
wire  wire175 = wire169 & wire174;
wire  wire176 = wire175 & wire63;
wire  wire177 = wire171 | wire176;
wire [7:0] wire178 = wire171 ? wire172 : wire65;
wire  wire179 = ~ wire63;
wire  wire180 = wire179 & wire123;
wire  wire181 = wire175 & wire180;
wire  wire182 = wire181 & wire71;
wire  wire183 = wire165 | wire182;
wire [7:0] wire184 = wire165 ? wire166 : wire38;
wire  wire185 = wire182 & wire74;
wire  wire186 = wire177 | wire185;
wire [7:0] wire187 = wire177 ? wire178 : wire76;
wire  wire188 = ~ wire74;
wire  wire189 = wire182 & wire188;
wire  wire190 = wire186 | wire189;
wire [7:0] wire191 = wire186 ? wire187 : wire12;
wire  wire192 = ~ wire71;
wire  wire193 = wire192 & wire121;
wire  wire194 = wire181 & wire193;
wire  wire195 = wire194 & wire82;
wire  wire196 = wire183 | wire195;
wire [7:0] wire197 = wire183 ? wire184 : wire38;
wire  wire198 = wire195 & wire86;
wire  wire199 = wire190 | wire198;
wire [7:0] wire200 = wire190 ? wire191 : wire88;
wire  wire201 = ~ wire86;
wire  wire202 = wire195 & wire201;
wire  wire203 = wire199 | wire202;
wire [7:0] wire204 = wire199 ? wire200 : wire12;
wire  wire205 = ~ wire82;
wire  wire206 = wire205 & wire119;
wire  wire207 = wire194 & wire206;
wire  wire208 = wire207 & wire94;
wire  wire209 = wire196 | wire208;
wire [7:0] wire210 = wire196 ? wire197 : wire38;
wire  wire211 = wire208 & wire99;
wire  wire212 = wire203 | wire211;
wire [7:0] wire213 = wire203 ? wire204 : wire101;
wire  wire214 = ~ wire99;
wire  wire215 = wire208 & wire214;
wire  wire216 = wire212 | wire215;
wire [7:0] wire217 = wire212 ? wire213 : wire12;
wire  wire218 = ~ wire94;
wire  wire219 = wire218 & wire117;
wire  wire220 = wire207 & wire219;
wire  wire221 = wire220 & wire107;
wire  wire222 = wire209 | wire221;
wire [7:0] wire223 = wire209 ? wire210 : wire38;
wire  wire224 = wire221 & wire110;
wire  wire225 = wire216 | wire224;
wire [7:0] wire226 = wire216 ? wire217 : wire112;
wire  wire227 = ~ wire110;
wire  wire228 = wire221 & wire227;
wire  wire229 = wire225 | wire228;
wire [7:0] wire230 = wire225 ? wire226 : wire12;
// effects 
assign guard = wire136;
assign value = wire0;
always@(posedge clk)
begin
	if(rst_n)
		begin
// reset 
		end
	else
		begin
	if(wire136)
		begin
// put  debug code here (display, stop, ...)
if(wire146) reg_4[wire29] <= wire28;
if(wire222) reg_3 <= wire223;
if(wire162) reg_2[wire163] <= wire164;
if(wire229) reg_1 <= wire230;
		end
		end
end
endmodule
